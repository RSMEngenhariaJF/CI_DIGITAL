module mapeia ();

    task ativa_saida (input [2:0]entrada, output [7:0]saida);
            assign saida = 8'b1;
    endtask

    
endmodule
module ieee754_adder_tb;
    reg [31:0] a, b,am,bm;
    wire [31:0] result,result_sub;
    wire [31:0] result_mult;
    ieee754_adder uut (
        .a(a),
        .b(b),
        .result(result)
    );

    ieee754_sub DUT(
    .a(a),
    .b(b),
    .result(result_sub)
    );

    ieee754_mult DUT2(
    .a(am),
    .b(bm),
    .result(result_mult)
    );

    initial begin
        // Teste de soma: 4,75 + 2,125 = 6,875 => 0_10000001_10111000000000000000000
        a = 32'b0_10000001_00110000000000000000000; // 4,75
        b = 32'b0_10000000_00010000000000000000000; // 2,125
        am = 32'b0_10000001_00110000000000000000000; // 4,75
        bm = 32'b0_10000000_00010000000000000000000; // 2,125
        //add_sub = 0; // Soma
        #10;
        $display("Soma: --> Sinal: %b -- Expoente: %b ---- Mantissa: %b", result[31], result[30:23], result[22:0]);

        // Teste de soma: 9,5 + 3,75 = 13,25 => 0_10000010_10101000000000000000000
        a = 32'b0_10000010_00110000000000000000000; // 9,5
        b = 32'b0_10000000_11100000000000000000000; // 3,75
        am = 32'b1_10000010_00110000000000000000000; // -9,5
        bm = 32'b0_10000000_11100000000000000000000; // 3,75
        #10;
        $display("Soma: --> Sinal: %b -- Expoente: %b ---- Mantissa: %b", result[31], result[30:23], result[22:0]);

         // Teste de soma: 3,75 - 9,5   = - 5,75 => 0_10000010_10101000000000000000000
        b = 32'b0_10000010_00110000000000000000000; // 9,5
        a = 32'b0_10000000_11100000000000000000000; // 3,75
        bm = 32'b0_10000010_00110000000000000000000; // 9,5
        am = 32'b1_10000000_11100000000000000000000; // -3,75
        #10;
        $display("Soma: --> Sinal: %b -- Expoente: %b ---- Mantissa: %b", result[31], result[30:23], result[22:0]);

         // Teste de soma: 9,75 - 9,75   = 0 => 0_10000010_10101000000000000000000
        a = 32'b0_10000010_00110000000000000000000; // 9,75
        b = 32'b0_10000010_00110000000000000000000; // 9,75
        am = 32'b0_10000010_00110000000000000000000; // 9,75
        bm = 32'b0_00000000_00000000000000000000000; // 9,75
        #10;



        $display("Soma: --> Sinal: %b -- Expoente: %b ---- Mantissa: %b", result[31], result[30:23], result[22:0]);
        $stop;
    end
endmodule


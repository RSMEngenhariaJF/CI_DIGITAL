module myand(
        input a,b,
        output x
);

assign x = a & b; 

endmodule 

`timescale 1ns / 100ps
module tb_conv_GRAY();

reg [3:0] bcd;
wire [3:0] S;

conv_gray DUT(
    .bcd,
    .S
    );

initial begin
    bcd = 4'b0000;
    #10 bcd = 4'b0000;
    #10 bcd = 4'b0001;
    #10 bcd = 4'b0010;
    #10 bcd = 4'b0011;
    #10 bcd = 4'b0100;
    #10 bcd = 4'b0101;
    #10 bcd = 4'b0110;
    #10 bcd = 4'b0111;
    #10 bcd = 4'b1000;
    #10 bcd = 4'b1001;
    #10 bcd = 4'b1010;
    #10 bcd = 4'b1011;
    #10 bcd = 4'b1100;
    #10 bcd = 4'b1101;
    #10 bcd = 4'b1110;
    #10 bcd = 4'b1111;
    #10 bcd = 4'b1111;
    $stop();
end 

endmodule
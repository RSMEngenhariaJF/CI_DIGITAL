module inv(
output b,
input a
);

assign b = ~a;

endmodule
module carry_look_ahead_adder_param #(parameter N) (
        input [N-1:0] A, //! Entrada A (4 bits)
        input [N-1:0] B, //! Entrada B (4 bits)
        input C_in , //! Carry inicial
        output [N-1:0] S, //! Soma final (4 bits)
        output C_out //! Carry final
);
 // Sinais intermediários para Carry -Generate (G) e  Carry -Propagate (P)
 wire [N-1:0] G; //! Carry -Generate
 wire [N-1:0] P; //! Carry -Propagate
 wire [N:0] C; //! Carry intermediário (C[0] = C_in , C[4] = 
 
 // Associar o Carry de entrada
 assign C[0] = C_in;
// Calcular G e P
 assign G = A & B; // G_i = A_i AND B_i
 assign P = A | B; // P_i = A_i OR B_i

    genvar i;
    generate
        for (i = 0; i < N; i = i + 1) begin 
            assign C[i+1] = G[i] | (P[i] & C[i]);
        end
    endgenerate
 // Calcular a soma
 assign S = A ^ B ^ C[N-1:0]; // S_i = A_i XOR B_i XOR C_i

 // Associar o Carry final
 assign C_out = C[N];
 endmodule

 module subtrator #(parameter N=4)(
        input [N-1:0] A,B,
        input B_in,
        output [N-1:0] D,
        output B_out
 );
    wire [N-1:0] B_comp, Dif;
    wire B_int;
    assign B_comp = (~B) +1'b1;
    
    carry_look_ahead_adder_param #(N) soma (
        .A(A), //! Entrada A (4 bits)
        .B(B_comp), //! Entrada B (4 bits)
        .C_in(B_in) , //! Carry inicial
        .S(Dif), //! Soma final (4 bits)
        .C_out(B_int) //! Carry final
    );

    assign {B_out,D} = {~B_int,Dif}; 

 endmodule
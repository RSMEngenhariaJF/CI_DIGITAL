module myand(
        input a,b,
        output x
);

x = a & b; 

endmodule 
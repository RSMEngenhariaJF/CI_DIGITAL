module dec_4_16 (
    input [3:0] A,
    output [15:0] S
);

reg [15:0] saida;

always @ (*) begin
    case (A)
            4'b0000 : saida <= 16'b10000000_00000000;
            4'b0001 : saida <= 16'b01000000_00000000;
            4'b0010 : saida <= 16'b00100000_00000000;
            4'b0011 : saida <= 16'b00010000_00000000;
            4'b0100 : saida <= 16'b00001000_00000000;
            4'b0101 : saida <= 16'b00000100_00000000;
            4'b0110 : saida <= 16'b00000010_00000000;
            4'b0111 : saida <= 16'b00000001_00000000;
            4'b1000 : saida <= 16'b00000000_10000000;
            4'b1001 : saida <= 16'b00000000_01000000;
            4'b1010 : saida <= 16'b00000000_00100000;
            4'b1011 : saida <= 16'b00000000_00010000;
            4'b1100 : saida <= 16'b00000000_00001000;
            4'b1101 : saida <= 16'b00000000_00000100;
            4'b1110 : saida <= 16'b00000000_00000010;
            4'b1111 : saida <= 16'b00000000_00000001;
            default: saida <=  16'b00000000_00000000;
    endcase
end

assign S = saida;

endmodule
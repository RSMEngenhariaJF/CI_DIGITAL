module conv_7seg(
    input [3:0] bcd,
    output [6:0] S
    );
    reg [7:0] Y;
    always @(*) begin
        case (bcd)
                4'b0000 : Y <= 7'b0000001;
                4'b0001 : Y <= 7'b1001111;
                4'b0010 : Y <= 7'b0010010;
                4'b0011 : Y <= 7'b0000110;
                4'b0100 : Y <= 7'b1001100;
                4'b0101 : Y <= 7'b0100100;
                4'b0110 : Y <= 7'b0100000;
                4'b0111 : Y <= 7'b0001111;
                4'b1000 : Y <= 7'b0000000;
                4'b1001 : Y <= 7'b0000100;
                4'b1010 : Y <= 7'b1111;
                4'b1011 : Y <= 7'b1110;
                4'b1100 : Y <= 7'b1010;
                4'b1101 : Y <= 7'b1011;
                4'b1110 : Y <= 7'b1001;
                4'b1111 : Y <= 7'b1000;
                
                default: Y <= 4'b0000; 
        endcase 
    end
    assign S = Y;
endmodule